//dddd
module ();

endmodule
